module MiniLab0_tb ();
    
endmodule
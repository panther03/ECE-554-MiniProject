localparam DMEM_DEPTH = 13;
localparam IMEM_DEPTH = 14;